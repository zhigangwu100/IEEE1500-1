module WBR1 (resetn,CLK,WPSI1,wse_outputs,hold_outputs,CoreOut,WPSO1,Dout);
input resetn;
input CLK;
input WPSI1;
//input ScanEnable;
//input HoldEnable;
input wse_outputs;
input hold_outputs;
input [7:0]CoreOut;
output WPSO1;
output [7:0]Dout;
wire [6:0]WBR1_connect;
//WC_SF1_CII DIN0(resetn,CLK,CoreOut[0],WPSI1,          ScanEnable,HoldEnable,Dout[0],WBR1_connect[0]);
//WC_SF1_CII DIN1(resetn,CLK,CoreOut[1],WBR1_connect[0],ScanEnable,HoldEnable,Dout[1],WBR1_connect[1]);
//WC_SF1_CII DIN2(resetn,CLK,CoreOut[2],WBR1_connect[1],ScanEnable,HoldEnable,Dout[2],WBR1_connect[2]);
//WC_SF1_CII DIN3(resetn,CLK,CoreOut[3],WBR1_connect[2],ScanEnable,HoldEnable,Dout[3],WBR1_connect[3]);
//WC_SF1_CII DIN4(resetn,CLK,CoreOut[4],WBR1_connect[3],ScanEnable,HoldEnable,Dout[4],WBR1_connect[4]);
//WC_SF1_CII DIN5(resetn,CLK,CoreOut[5],WBR1_connect[4],ScanEnable,HoldEnable,Dout[5],WBR1_connect[5]);
//WC_SF1_CII DIN6(resetn,CLK,CoreOut[6],WBR1_connect[5],ScanEnable,HoldEnable,Dout[6],WBR1_connect[6]);
//WC_SF1_CII DIN7(resetn,CLK,CoreOut[7],WBR1_connect[6],ScanEnable,HoldEnable,Dout[7],WPSO1);
WC_SF1_CII DOUT0(resetn,CLK,CoreOut[0],WPSI1,          wse_outputs,hold_outputs,Dout[0],WBR1_connect[0]);
WC_SF1_CII DOUT1(resetn,CLK,CoreOut[1],WBR1_connect[0],wse_outputs,hold_outputs,Dout[1],WBR1_connect[1]);
WC_SF1_CII DOUT2(resetn,CLK,CoreOut[2],WBR1_connect[1],wse_outputs,hold_outputs,Dout[2],WBR1_connect[2]);
WC_SF1_CII DOUT3(resetn,CLK,CoreOut[3],WBR1_connect[2],wse_outputs,hold_outputs,Dout[3],WBR1_connect[3]);
WC_SF1_CII DOUT4(resetn,CLK,CoreOut[4],WBR1_connect[3],wse_outputs,hold_outputs,Dout[4],WBR1_connect[4]);
WC_SF1_CII DOUT5(resetn,CLK,CoreOut[5],WBR1_connect[4],wse_outputs,hold_outputs,Dout[5],WBR1_connect[5]);
WC_SF1_CII DOUT6(resetn,CLK,CoreOut[6],WBR1_connect[5],wse_outputs,hold_outputs,Dout[6],WBR1_connect[6]);
WC_SF1_CII DOUT7(resetn,CLK,CoreOut[7],WBR1_connect[6],wse_outputs,hold_outputs,Dout[7],WPSO1);
endmodule